//ALL_TIME
//controls all time related commands

module	ALL_TIME	(	
		input	logic	clk,
		input	logic	resetN,
		input	logic	run,      //game is running
		input logic turbo,    //sets the game to turbo mode
		input	logic	Ice,      //freeze enemy advancment and spawn
		
		output logic spawn,   //the rate of creation of new enemies
		output logic advance, //the speed of advancment
		output logic lvl      //current lvl of the game
);


//Fill your code here



endmodule
